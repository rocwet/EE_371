library verilog;
use verilog.vl_types.all;
entity ripple_down_vlg_check_tst is
    port(
        Q_0             : in     vl_logic;
        Q_1             : in     vl_logic;
        Q_2             : in     vl_logic;
        Q_3             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ripple_down_vlg_check_tst;
