library verilog;
use verilog.vl_types.all;
entity ripple_down_vlg_vec_tst is
end ripple_down_vlg_vec_tst;
