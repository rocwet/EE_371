library verilog;
use verilog.vl_types.all;
entity johnson_down_vlg_vec_tst is
end johnson_down_vlg_vec_tst;
