module test(out, in1);
	output out;
	input in1;
	
	assign out = in1;



endmodule 